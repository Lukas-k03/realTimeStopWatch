module finalOutput();

endmodule